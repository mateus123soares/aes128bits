library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity shiftRows is
	
	 port(
		mensagem: in std_logic_vector(127 downto 0); --mensagem a ser codificada
		saida: out std_logic_vector(127 downto 0)	--saida
		);

end shiftRows;

architecture Behavior of shiftRows is
	
	signal shift,shift2,shift3,shift4: std_logic_vector(31 downto 0);
	signal palavra,palavra2,palavra3,palavra4: std_logic_vector(31 downto 0);
	
	begin
	
	shift <= mensagem(127 downto 96);
	shift2 <= mensagem(95 downto 64);
	shift3 <= mensagem(63 downto 32);
	shift4 <= mensagem(31 downto 0);
	
	palavra <= shift(31 downto 24) & shift2(23 downto 16) & shift3(15 downto 8) & shift4(7 downto 0);
	palavra2 <= shift2(31 downto 24) & shift3(23 downto 16) & shift4(15 downto 8) & shift(7 downto 0);
	palavra3 <= shift3(31 downto 24) & shift4(23 downto 16) & shift(15 downto 8) & shift2(7 downto 0);
	palavra4 <= shift4(31 downto 24) & shift(23 downto 16) & shift2(15 downto 8)  & shift3(7 downto 0);
	
	saida <= palavra & palavra2 & palavra3 & palavra4;
	
end Behavior;
	